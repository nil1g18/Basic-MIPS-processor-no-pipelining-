`define N_BIT 16
`define PC_SIZE 16
`define INSTR_SIZE 32
`define PC_INCREMENT 1

`define ALU_FUNC_SIZE 3

`define REG_ADDR_SIZE 6

`define REG_ZERO 0